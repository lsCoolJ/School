library verilog;
use verilog.vl_types.all;
entity testLaser16 is
end testLaser16;

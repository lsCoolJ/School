library verilog;
use verilog.vl_types.all;
entity testCountdownTimer is
end testCountdownTimer;

library verilog;
use verilog.vl_types.all;
entity Test_Mux3w5to1 is
end Test_Mux3w5to1;

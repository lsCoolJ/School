library verilog;
use verilog.vl_types.all;
entity testBCDAdd is
end testBCDAdd;

library verilog;
use verilog.vl_types.all;
entity testCountNG is
end testCountNG;

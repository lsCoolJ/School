/*Homework 1 Part 2 by Ben Foster
 *TCES 330 4/16/14
 */
module HW1Part2(SW, LEDR, LEDG);
	input [17:0] SW; //Toggle switches
	output [17:0] LEDR; //Red LEDs
	output [7:0] LEDG; //Green LEDs
	wire S; //Select line
	
	assign S = SW[17]; //assign select line to last switch
	assign LEDR = SW; //know which switch is on
	
	//Instance of the Mux
	Mux8 I1(S, SW[7:0], SW[15:8], LEDG[7:0]);
	
endmodule

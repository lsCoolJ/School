//------------------------------------------------------------------
//
// TCES 330, Spring 2011
// R. Gutmann
// 
// This module is the testbench for RegisterFile
// Used in our processor, tested with ModelSim
//
//------------------------------------------------------------------

`timescale 1 ns/1 ns
module testRegisterFile();
	
	//DUT inputs:
	reg Clk;		// system clock;
	reg Rst;		// register file reset (everything to zero)
	reg Wen;		// write enable (enable write side decoder)
	reg [3:0] WAddr;	//write address (which register to write to)
	reg [15:0] WData;	// data to write to a register
	reg [3:0] RAAddr, RBAddr;	// which regisers to read from
	reg RAen, RBen;				// A and B-side read enables
	
	//DUT outputs
	wire [15:0] RAData, RBData;	//A- and B-side read data
	
	//reference RegisterFile( Clk, Rst, W_en, W_Addr, W_Data, Ra_Addr, Rb_Addr, Ra_en, Ra_Data, Rb_Data);
	RegisterFile DUT( Clk, Rst, Wen, WAddr, WData, RAAddr, RBAddr, RAen, RBen, RAData, RBData );
	
	// generate clock
	always begin
		Clk = 0;
		#10;
		Clk = 1'b1;
		#10;
	end
	
	integer I;
	
	initial begin
		//load up the registers
		Rst = 1;
		#20 Rst = 0;
		#20 for (I = 0; I < 16; I = I + 1) begin
			#20 WData = I + 16'h10;
			WAddr = I;
			Wen = 1;
			#20 Wen = 0;
		end
		
		//read the registers
		#20 for(I = 0; I < 16; I = I + 1) begin
			#20 RAAddr = I;
			RBAddr = (I + 4'h8) % 16;
			RAen = 1;
			RBen = 1;
			#20 RAen = 0;
			RBen = 0;
		end
		#20 $stop;
	end //initial
	
endmodule

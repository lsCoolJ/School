library verilog;
use verilog.vl_types.all;
entity testDragRace is
end testDragRace;

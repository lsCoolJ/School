library verilog;
use verilog.vl_types.all;
entity testALU is
end testALU;

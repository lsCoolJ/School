library verilog;
use verilog.vl_types.all;
entity testMux5 is
end testMux5;

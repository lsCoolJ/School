library verilog;
use verilog.vl_types.all;
entity testRegisterFile is
end testRegisterFile;
